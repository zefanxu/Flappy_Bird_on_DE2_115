//-------------------------------------------------------------------------
//    Color_Mapper.sv                                                    --
//    Stephen Kempf                                                      --
//    3-1-06                                                             --
//                                                                       --
//    Modified by David Kesler  07-16-2008                               --
//    Translated by Joe Meng    07-07-2013                               --
//                                                                       --
//    Fall 2014 Distribution                                             --
//                                                                       --
//    For use with ECE 385 Lab 7                                         --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------

    
module  color_mapper ( input        [9:0] PipePositionX, PipePositionY, DrawX, DrawY, Ball_size,
                       output logic [7:0]  Red, Green, Blue );
    
    logic pipe_green_on;
	 
 /* Old Ball: Generated square box by checking if the current pixel is within a square of length
    2*Ball_Size, centered at (BallX, BallY).  Note that this requires unsigned comparisons.
	 
    if ((DrawX >= BallX - Ball_size) &&
       (DrawX <= BallX + Ball_size) &&
       (DrawY >= BallY - Ball_size) &&
       (DrawY <= BallY + Ball_size))

     New Ball: Generates (pixelated) circle by using the standard circle formula.  Note that while 
     this single line is quite powerful descriptively, it causes the synthesis tool to use up three
     of the 12 available multipliers on the chip!  Since the multiplicants are required to be signed,
	  we have to first cast them from logic to int (signed by default) before they are multiplied). */
	  
    

	PipesGreenBodyTop <= (DrawX>=PipePositionX+12) && (DrawX<=PipePositionX+78) && (DrawY>=0) && (DrawY<=PipePositionY);
    PipesGreenTop <= (CounterX>=PipePositionX+3) && (CounterX<=PipePositionX+87) && (CounterY>=PipePositionY+3) && (CounterY<=PipePositionY+30);

    always_comb
    begin:pipe_green_on_proc
        if ( PipesGreenTop || PipesGreenBodyTop ) 
            pipe_green_on = 1'b1;
        else 
            pipe_green_on = 1'b0;
     end 
       
    always_comb
    begin:RGB_Display
        if ((pipe_green_on == 1'b1)) 
        begin 
            Red = 8'h00;
            Green = 8'hff;
            Blue = 8'h00;
        end       
        else 
        begin 
            Red = 8'h3f; 
            Green = 8'h00;
            Blue = 8'h3f - DrawX[9:3];
        end      
    end 
    
endmodule
